module Tail_light (CLK,RST,LEFT,RIGHT,HAZ,LA,LB,LC,RA,RB,RC ) ;
input CLK,RST,LEFT,RIGHT,HAZ;
output reg LA,LB,LC,RA,RB, RC;
reg[2:0]Sreg,Snext;

parameter [2:0]IDLE=3'b000,L1=3'b001,L2=3'b011,L3=3'b010,
					R1=3'b101,R2=3'b111,R3=3'b110,LR3=3'b100;
wire CLK_1HzOut;
Divider50MHz uD50(CLK, RST, CLK_1HzOut);
always@(posedge CLK_1HzOut or negedge RST)//时序逻辑:存储状态
begin
if(~RST)Sreg <= IDLE;
else Sreg <= Snext;
end
always@ (LEFT,RIGHT,HAZ,Sreg)begin
case(Sreg)IDLE:if(HAZ|(LEFT&RIGHT))Snext=LR3;
			else if(RIGHT)Snext= R1;
			else if(LEFT)Snext= L1;
			else Snext = IDLE;
			R1:Snext= R2;
			R2:Snext= R3;
			R3:Snext= IDLE;
			L1:Snext =L2;
			L2:Snext= L3;
				L3:Snext= IDLE;
			LR3:Snext= IDLE;
			default:Snext = IDLE;
endcase
end
always @(Sreg)begin
case(Sreg)
IDLE:{LC,LB,LA,RA,RB,RC}= 6'b00_0000;
R1:{LC,LB,LA,RA,RB,RC}= 6'b00_0100;
R2:{LC,LB,LA,RA,RB,RC}= 6'b00_0110;
R3:{LC,LB,LA,RA,RB,RC}= 6'b00_0111;
L1:{LC,LB,LA,RA,RB,RC}= 6'b00_1000;
L2:{LC,LB,LA,RA,RB,RC}= 6'b01_1000;
L3:{LC,LB,LA,RA,RB,RC}= 6'b11_1000;
LR3:{LC,LB,LA,RA,RB,RC}= 6'b11_1111;
default:{LC,LB,LA,RA,RB,RC}=6'b00_0000;
endcase
end
endmodule
